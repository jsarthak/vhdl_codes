LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY nor_gate IS
    PORT (
        a, b : IN STD_LOGIC;
        y : OUT STD_LOGIC);
END nor_gate;

ARCHITECTURE DataFlow OF nor_gate IS

BEGIN

    y <= a NOR b;

END DataFlow;