LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY xor_gate IS
    PORT (
        a, b : IN STD_LOGIC;
        y : OUT STD_LOGIC);
END xor_gate;

ARCHITECTURE Behavioral OF xor_gate IS

BEGIN
    y <= a XOR b;

END Behavioral;