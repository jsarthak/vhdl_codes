LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ex3 IS
    PORT (
        BCD : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        EXCESS : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END ex3;

ARCHITECTURE Behavioral OF ex3 IS
BEGIN
    PROCESS (BCD)
    BEGIN
        IF (BCD > "1001") THEN
            EXCESS <= "XXXX";
        ELSE
            EXCESS <= BCD + 3;
        END IF;
    END PROCESS;
END Behavioral;